VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO power_switch
  CLASS BLOCK ;
  FOREIGN power_switch ;
  ORIGIN 12.120 37.580 ;
  SIZE 43.250 BY 53.870 ;
  PIN gate
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -2.570 0.360 -2.270 11.300 ;
    END
  END gate
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -12.120 -37.580 -5.560 15.860 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.560 -37.220 31.130 16.290 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT -0.085 -0.085 17.025 11.745 ;
      LAYER met1 ;
        RECT -2.270 11.580 20.120 12.000 ;
        RECT -1.990 0.080 20.120 11.580 ;
        RECT -2.270 -0.190 20.120 0.080 ;
      LAYER met2 ;
        RECT -1.090 -1.970 17.830 14.470 ;
      LAYER met3 ;
        RECT -1.020 -2.900 17.630 14.460 ;
      LAYER met4 ;
        RECT -5.160 -6.280 23.160 16.180 ;
  END
END power_switch
END LIBRARY

