magic
tech sky130A
magscale 1 2
timestamp 1684691938
<< metal1 >>
rect 82 2368 3308 2372
rect 3636 2368 4024 2400
rect 82 2366 4024 2368
rect 54 2294 60 2366
rect 3338 2340 4024 2366
rect 3338 2308 3696 2340
rect 3338 2294 3344 2308
rect -514 2200 3310 2260
rect -514 132 -454 2200
rect -218 2052 3562 2132
rect -218 1402 -128 2052
rect 3472 1402 3562 2052
rect -218 1270 3562 1402
rect -214 940 3566 1066
rect -214 290 -122 940
rect 3478 290 3566 940
rect -214 204 3566 290
rect -514 130 154 132
rect -514 72 3312 130
rect 86 70 3312 72
rect 3964 22 4024 2340
rect 86 -38 4024 22
<< via1 >>
rect 60 2294 3338 2366
rect -128 1402 3472 2052
rect -122 290 3478 940
<< metal2 >>
rect -192 2366 3540 2894
rect -192 2294 60 2366
rect 3338 2294 3540 2366
rect -192 2132 3540 2294
rect -218 2052 3562 2132
rect -218 1402 -128 2052
rect 3472 1402 3562 2052
rect -218 1270 3562 1402
rect -214 940 3566 1066
rect -214 290 -122 940
rect 3478 290 3566 940
rect -214 204 3566 290
rect -206 -394 3526 204
use sky130_fd_pr__pfet_01v8_7HKEJJ  sky130_fd_pr__pfet_01v8_7HKEJJ_0
timestamp 1684691938
transform 1 0 1694 0 1 1166
box -1747 -1219 1747 1219
<< labels >>
flabel metal2 -192 2052 3540 2894 0 FreeSans 800 0 0 0 source
port 0 nsew
flabel metal2 -206 -394 3526 290 0 FreeSans 800 0 0 0 drain
port 1 nsew
flabel metal1 -514 72 -454 2260 0 FreeSans 800 0 0 0 gate
port 2 nsew
<< end >>
